//
//  configurations
//
//
`define RESET_VECTOR        'h00000000

//
//  instruction patterns
//
//
`define INST_PATTERN_LUI    'b?????????????????????????0110111

`define INST_PATTERN_AUIPC  'b?????????????????????????0010111

`define INST_PATTERN_JAL    'b?????????????????????????1101111

`define INST_PATTERN_JALR   'b?????????????????000?????1100111

`define INST_PATTERN_BRANCH 'b?????????????????????????1100011
`define INST_PATTERN_BEQ    'b?????????????????000?????1100011
`define INST_PATTERN_BNE    'b?????????????????001?????1100011
`define INST_PATTERN_BLT    'b?????????????????100?????1100011
`define INST_PATTERN_BGE    'b?????????????????101?????1100011
`define INST_PATTERN_BLTU   'b?????????????????110?????1100011
`define INST_PATTERN_BGEU   'b?????????????????111?????1100011

`define INST_PATTERN_LOAD   'b?????????????????????????0000011
`define INST_PATTERN_LB     'b?????????????????000?????0000011
`define INST_PATTERN_LH     'b?????????????????001?????0000011
`define INST_PATTERN_LW     'b?????????????????010?????0000011
`define INST_PATTERN_LBU    'b?????????????????100?????0000011
`define INST_PATTERN_LHU    'b?????????????????101?????0000011

`define INST_PATTERN_STORE  'b?????????????????????????0100011
`define INST_PATTERN_SB     'b?????????????????000?????0100011
`define INST_PATTERN_SH     'b?????????????????001?????0100011
`define INST_PATTERN_SW     'b?????????????????010?????0100011

`define INST_PATTERN_ALGI   'b?????????????????????????0010011
`define INST_PATTERN_ADDI   'b?????????????????000?????0010011
`define INST_PATTERN_SLTI   'b?????????????????010?????0010011
`define INST_PATTERN_SLTIU  'b?????????????????011?????0010011
`define INST_PATTERN_XORI   'b?????????????????100?????0010011
`define INST_PATTERN_ORI    'b?????????????????110?????0010011
`define INST_PATTERN_ANDI   'b?????????????????111?????0010011
`define INST_PATTERN_SLLI   'b0000000??????????001?????0010011
`define INST_PATTERN_SRLI   'b0000000??????????101?????0010011
`define INST_PATTERN_SRAI   'b0100000??????????101?????0010011

`define INST_PATTERN_ALG    'b?????????????????????????0110011
`define INST_PATTERN_ADD    'b0000000??????????000?????0110011
`define INST_PATTERN_SUB    'b0100000??????????000?????0110011
`define INST_PATTERN_SLL    'b0000000??????????001?????0110011
`define INST_PATTERN_SLT    'b0000000??????????010?????0110011
`define INST_PATTERN_SLTU   'b0000000??????????011?????0110011
`define INST_PATTERN_XOR    'b0000000??????????100?????0110011
`define INST_PATTERN_SRL    'b0000000??????????101?????0110011
`define INST_PATTERN_SRA    'b0100000??????????101?????0110011
`define INST_PATTERN_OR     'b0000000??????????110?????0110011
`define INST_PATTERN_AND    'b0000000??????????111?????0110011

`define INST_PATTERN_SYNCH  'b?????????????????????????0001111
`define INST_PATTERN_FENCE  'b0000????????00000000000000001111
`define INST_PATTERN_FENCEI 'b00000000000000000001000000001111

`define INST_PATTERN_SYSTEM 'b?????????????????????????1110011
`define INST_PATTERN_ECALL  'b00000000000000000000000001110011
`define INST_PATTERN_EBREAK 'b00000000000100000000000001110011
`define INST_PATTERN_CSRRW  'b?????????????????001?????1110011
`define INST_PATTERN_CSRRS  'b?????????????????010?????1110011
`define INST_PATTERN_CSRRC  'b?????????????????011?????1110011
`define INST_PATTERN_CSRRWI 'b?????????????????101?????1110011
`define INST_PATTERN_CSRRSI 'b?????????????????110?????1110011
`define INST_PATTERN_CSRRCI 'b?????????????????111?????1110011

