`define ALU_OP_ADD  'b0000
`define ALU_OP_SUB  'b1000
`define ALU_OP_SLL  'b0001
`define ALU_OP_SLT  'b0010
`define ALU_OP_SLTU 'b0011
`define ALU_OP_XOR  'b0100
`define ALU_OP_SRL  'b0101
`define ALU_OP_SRA  'b1101
`define ALU_OP_OR   'b0110
`define ALU_OP_AND  'b0111

`define BALU_OP_EQ  'b000
`define BALU_OP_NE  'b001
`define BALU_OP_LT  'b100
`define BALU_OP_GE  'b101
`define BALU_OP_LTU 'b110
`define BALU_OP_GEU 'b111

